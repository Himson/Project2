`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/22/2019 03:51:05 PM
// Design Name: 
// Module Name: mux2to1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux2to1(
    input [31:0] port0,
    input [31:0] port1,
    input control,
    output reg[31:0] out 
    );
    always@(*)begin
        case(control)
            1'b0: out = port0;
            1'b1: out = port1;
            default: out = port0;
        endcase
    end
endmodule
